`include "comm_param.svh"

`include "comm_param.vh"

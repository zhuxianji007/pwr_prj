`include "com_param.svh"

parameter LV_SCAN_REG_NUM           = 6                                                         ,

parameter EFUSE_DATA_NUM            = 8                                                         ,
parameter EFUSE_DW                  = REG_DW                                                    ,

parameter HV_ANALOG_REG_START_ADDR  = 7'h40                                                     ,
parameter HV_ANALOG_REG_END_ADDR    = 7'h6E                                                     ,

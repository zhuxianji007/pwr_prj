//============================================================
//Module   : lv_pkg
//Function : define structure
//File Tree: 
//-------------------------------------------------------------
//Update History
//-------------------------------------------------------------
//Rev.level     Date          Code_by         Contents
//1.0           2022/11/6     xxxx            Create
//=============================================================

`ifndef LV_PKG_SV
`defien LV_PKG_SV

package lv_pkg;

    import com_pkg::*;

endpackage

`endif //LV_PKG_SV

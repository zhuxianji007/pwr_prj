`include "comm_param.svh"

parameter EFUSE_DATA_NUM        = 16                                                        ,
parameter EFUSE_DW              = REG_DW                                                    ,

sxx
